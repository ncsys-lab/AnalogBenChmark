

module comparator_latch #
(
  parameter n_to_response_time = -1038,
  parameter p_to_response_time = -1020,
  parameter const_response_time = 1285,
  parameter n_to_tau = -1248,
  parameter p_to_tau = 1037,
  parameter const_tau = 1042,
  parameter n_to_response_time_lh = -1752,
  parameter p_to_response_time_lh = -1006,
  parameter const_response_time_lh = 1185,
  parameter n_to_tau_lh = 1131,
  parameter p_to_tau_lh = -1115,
  parameter const_tau_lh = 1529
)
(
  input clk,
  input reset,
  input sys_clk,
  input [10-1:0] n,
  input [10-1:0] p,
  output [10-1:0] out
);

  reg [17-1:0] state_cycle_counter;
  reg [1-1:0] prev_sys_clk;
  reg [35-1:0] o;
  wire [32-1:0] wait_time;
  wire [51-1:0] tau;
  wire [36-1:0] dvdt;
  wire [32-1:0] wait_time_lh;
  wire [59-1:0] tau_lh;
  wire [37-1:0] dodt;
  reg [32-1:0] fsm;
  localparam fsm_init = 0;
  wire [35-1:0] padr_0;
  wire [20-1:0] padr_bits_1;
  assign padr_bits_1 = 0;
  wire [43-1:0] truncR_2;
  wire [43-1:0] padl_3;
  wire [41-1:0] padl_bits_4;
  wire [1-1:0] toSInt_5;
  assign toSInt_5 = 0;
  wire [41-1:0] toSInt_imm_6;
  wire [40-1:0] const_7;
  assign const_7 = 40'd907097092915;
  assign toSInt_imm_6 = { toSInt_5, const_7 };
  assign padl_bits_4 = toSInt_imm_6;
  assign padl_3 = { { 2{ padl_bits_4[40] } }, padl_bits_4 };
  assign truncR_2 = padl_3;
  wire [15-1:0] truncR_shift_8;
  assign truncR_shift_8 = truncR_2 >>> 28;
  wire [15-1:0] truncR_imm_9;
  assign truncR_imm_9 = (truncR_2[42])? truncR_shift_8[14:0] : truncR_2[42:28];
  assign padr_0 = { truncR_imm_9, padr_bits_1 };
  wire [13-1:0] truncR_10;
  wire [14-1:0] truncval_11;
  wire [15-1:0] toUsInt_12;
  wire [35-1:0] truncR_13;
  assign truncR_13 = o;
  wire [15-1:0] truncR_shift_14;
  assign truncR_shift_14 = truncR_13 >>> 20;
  wire [15-1:0] truncR_imm_15;
  assign truncR_imm_15 = (truncR_13[34])? truncR_shift_14[14:0] : truncR_13[34:20];
  assign toUsInt_12 = truncR_imm_15;
  assign truncval_11 = toUsInt_12[11:0];
  assign truncR_10 = truncval_11[12:0];
  wire [32-1:0] padl_16;
  wire [18-1:0] padl_bits_17;
  wire [39-1:0] truncR_18;
  wire [39-1:0] padl_19;
  wire [24-1:0] padl_bits_20;
  wire [117-1:0] truncR_21;
  wire [184-1:0] truncval_22;
  wire [184-1:0] padl_23;
  wire [92-1:0] padl_bits_24;
  wire [92-1:0] padl_25;
  wire [59-1:0] padl_bits_26;
  wire [98-1:0] truncR_27;
  wire [105-1:0] truncval_28;
  wire [105-1:0] padl_29;
  wire [52-1:0] padl_bits_30;
  wire [52-1:0] padr_31;
  wire [41-1:0] padr_bits_32;
  assign padr_bits_32 = 0;
  wire [1-1:0] toSInt_33;
  assign toSInt_33 = 0;
  wire [11-1:0] toSInt_imm_34;
  assign toSInt_imm_34 = { toSInt_33, n };
  assign padr_31 = { toSInt_imm_34, padr_bits_32 };
  assign padl_bits_30 = padr_31;
  assign padl_29 = { { 53{ padl_bits_30[51] } }, padl_bits_30 };
  wire [105-1:0] padl_35;
  wire [52-1:0] padl_bits_36;
  wire [52-1:0] padl_37;
  wire [50-1:0] padl_bits_38;
  wire [50-1:0] param_39;
  assign param_39 = n_to_response_time;
  assign padl_bits_38 = param_39;
  assign padl_37 = { { 2{ padl_bits_38[49] } }, padl_bits_38 };
  assign padl_bits_36 = padl_37;
  assign padl_35 = { { 53{ padl_bits_36[51] } }, padl_bits_36 };
  assign truncval_28 = padl_29 * padl_35;
  wire [98-1:0] truncval_imm_40;
  assign truncval_imm_40 = { truncval_28[104], truncval_28[96:0] };
  assign truncR_27 = truncval_imm_40;
  wire [59-1:0] truncR_shift_41;
  assign truncR_shift_41 = truncR_27 >>> 39;
  wire [59-1:0] truncR_imm_42;
  assign truncR_imm_42 = (truncR_27[97])? truncR_shift_41[58:0] : truncR_27[97:39];
  wire [59-1:0] padr_43;
  wire [2-1:0] padr_bits_44;
  assign padr_bits_44 = 0;
  wire [94-1:0] truncR_45;
  wire [101-1:0] truncval_46;
  wire [101-1:0] padl_47;
  wire [50-1:0] padl_bits_48;
  wire [50-1:0] padr_49;
  wire [39-1:0] padr_bits_50;
  assign padr_bits_50 = 0;
  wire [1-1:0] toSInt_51;
  assign toSInt_51 = 0;
  wire [11-1:0] toSInt_imm_52;
  assign toSInt_imm_52 = { toSInt_51, p };
  assign padr_49 = { toSInt_imm_52, padr_bits_50 };
  assign padl_bits_48 = padr_49;
  assign padl_47 = { { 51{ padl_bits_48[49] } }, padl_bits_48 };
  wire [101-1:0] padl_53;
  wire [50-1:0] padl_bits_54;
  wire [50-1:0] padl_55;
  wire [48-1:0] padl_bits_56;
  wire [48-1:0] param_57;
  assign param_57 = p_to_response_time;
  assign padl_bits_56 = param_57;
  assign padl_55 = { { 2{ padl_bits_56[47] } }, padl_bits_56 };
  assign padl_bits_54 = padl_55;
  assign padl_53 = { { 51{ padl_bits_54[49] } }, padl_bits_54 };
  assign truncval_46 = padl_47 * padl_53;
  wire [94-1:0] truncval_imm_58;
  assign truncval_imm_58 = { truncval_46[100], truncval_46[92:0] };
  assign truncR_45 = truncval_imm_58;
  wire [57-1:0] truncR_shift_59;
  assign truncR_shift_59 = truncR_45 >>> 37;
  wire [57-1:0] truncR_imm_60;
  assign truncR_imm_60 = (truncR_45[93])? truncR_shift_59[56:0] : truncR_45[93:37];
  assign padr_43 = { truncR_imm_60, padr_bits_44 };
  wire [59-1:0] padr_61;
  wire [15-1:0] padr_bits_62;
  assign padr_bits_62 = 0;
  wire [44-1:0] padl_63;
  wire [43-1:0] padl_bits_64;
  wire [1-1:0] toSInt_65;
  assign toSInt_65 = 0;
  wire [43-1:0] toSInt_imm_66;
  wire [42-1:0] param_67;
  assign param_67 = const_response_time;
  assign toSInt_imm_66 = { toSInt_65, param_67 };
  assign padl_bits_64 = toSInt_imm_66;
  assign padl_63 = { { 1{ padl_bits_64[42] } }, padl_bits_64 };
  assign padr_61 = { padl_63, padr_bits_62 };
  assign padl_bits_26 = truncR_imm_42 + padr_43 + padr_61;
  assign padl_25 = { { 33{ padl_bits_26[58] } }, padl_bits_26 };
  assign padl_bits_24 = padl_25;
  assign padl_23 = { { 92{ padl_bits_24[91] } }, padl_bits_24 };
  wire [184-1:0] padl_68;
  wire [92-1:0] padl_bits_69;
  wire [92-1:0] padr_70;
  wire [51-1:0] padr_bits_71;
  assign padr_bits_71 = 0;
  wire [1-1:0] toSInt_72;
  assign toSInt_72 = 0;
  wire [41-1:0] toSInt_imm_73;
  wire [40-1:0] const_74;
  assign const_74 = 40'd640000000000;
  assign toSInt_imm_73 = { toSInt_72, const_74 };
  assign padr_70 = { toSInt_imm_73, padr_bits_71 };
  assign padl_bits_69 = padr_70;
  assign padl_68 = { { 92{ padl_bits_69[91] } }, padl_bits_69 };
  assign truncval_22 = padl_23 * padl_68;
  assign truncR_21 = truncval_22[116:0];
  assign padl_bits_20 = truncR_21[116:93];
  wire [15-1:0] padl_bits_zero_75;
  assign padl_bits_zero_75 = 0;
  assign padl_19 = { padl_bits_zero_75, padl_bits_20 };
  assign truncR_18 = padl_19;
  assign padl_bits_17 = truncR_18[38:21];
  wire [14-1:0] padl_bits_zero_76;
  assign padl_bits_zero_76 = 0;
  assign padl_16 = { padl_bits_zero_76, padl_bits_17 };
  assign wait_time = padl_16;
  wire [35-1:0] padr_77;
  wire [20-1:0] padr_bits_78;
  assign padr_bits_78 = 0;
  wire [43-1:0] truncR_79;
  wire [43-1:0] padl_80;
  wire [41-1:0] padl_bits_81;
  wire [1-1:0] toSInt_82;
  assign toSInt_82 = 0;
  wire [41-1:0] toSInt_imm_83;
  wire [40-1:0] const_84;
  assign const_84 = 40'd907097092915;
  assign toSInt_imm_83 = { toSInt_82, const_84 };
  assign padl_bits_81 = toSInt_imm_83;
  assign padl_80 = { { 2{ padl_bits_81[40] } }, padl_bits_81 };
  assign truncR_79 = padl_80;
  wire [15-1:0] truncR_shift_85;
  assign truncR_shift_85 = truncR_79 >>> 28;
  wire [15-1:0] truncR_imm_86;
  assign truncR_imm_86 = (truncR_79[42])? truncR_shift_85[14:0] : truncR_79[42:28];
  assign padr_77 = { truncR_imm_86, padr_bits_78 };
  wire [13-1:0] truncR_87;
  wire [14-1:0] truncval_88;
  wire [15-1:0] toUsInt_89;
  wire [35-1:0] truncR_90;
  assign truncR_90 = o;
  wire [15-1:0] truncR_shift_91;
  assign truncR_shift_91 = truncR_90 >>> 20;
  wire [15-1:0] truncR_imm_92;
  assign truncR_imm_92 = (truncR_90[34])? truncR_shift_91[14:0] : truncR_90[34:20];
  assign toUsInt_89 = truncR_imm_92;
  assign truncval_88 = toUsInt_89[11:0];
  assign truncR_87 = truncval_88[12:0];
  wire [52-1:0] truncR_93;
  wire [53-1:0] truncval_94;
  wire [54-1:0] toUsInt_95;
  wire [54-1:0] padr_96;
  wire [1-1:0] padr_bits_97;
  assign padr_bits_97 = 0;
  wire [88-1:0] truncR_98;
  wire [95-1:0] truncval_99;
  wire [95-1:0] padl_100;
  wire [47-1:0] padl_bits_101;
  wire [47-1:0] padr_102;
  wire [36-1:0] padr_bits_103;
  assign padr_bits_103 = 0;
  wire [1-1:0] toSInt_104;
  assign toSInt_104 = 0;
  wire [11-1:0] toSInt_imm_105;
  assign toSInt_imm_105 = { toSInt_104, n };
  assign padr_102 = { toSInt_imm_105, padr_bits_103 };
  assign padl_bits_101 = padr_102;
  assign padl_100 = { { 48{ padl_bits_101[46] } }, padl_bits_101 };
  wire [95-1:0] padl_106;
  wire [47-1:0] padl_bits_107;
  wire [47-1:0] padl_108;
  wire [45-1:0] padl_bits_109;
  wire [45-1:0] param_110;
  assign param_110 = n_to_tau;
  assign padl_bits_109 = param_110;
  assign padl_108 = { { 2{ padl_bits_109[44] } }, padl_bits_109 };
  assign padl_bits_107 = padl_108;
  assign padl_106 = { { 48{ padl_bits_107[46] } }, padl_bits_107 };
  assign truncval_99 = padl_100 * padl_106;
  wire [88-1:0] truncval_imm_111;
  assign truncval_imm_111 = { truncval_99[94], truncval_99[86:0] };
  assign truncR_98 = truncval_imm_111;
  wire [53-1:0] truncR_shift_112;
  assign truncR_shift_112 = truncR_98 >>> 35;
  wire [53-1:0] truncR_imm_113;
  assign truncR_imm_113 = (truncR_98[87])? truncR_shift_112[52:0] : truncR_98[87:35];
  assign padr_96 = { truncR_imm_113, padr_bits_97 };
  wire [54-1:0] padl_114;
  wire [53-1:0] padl_bits_115;
  wire [1-1:0] toSInt_116;
  assign toSInt_116 = 0;
  wire [53-1:0] toSInt_imm_117;
  wire [86-1:0] truncR_118;
  wire [92-1:0] truncval_119;
  wire [92-1:0] padl_120;
  wire [46-1:0] padl_bits_121;
  wire [46-1:0] padr_122;
  wire [36-1:0] padr_bits_123;
  assign padr_bits_123 = 0;
  assign padr_122 = { p, padr_bits_123 };
  assign padl_bits_121 = padr_122;
  wire [46-1:0] padl_bits_zero_124;
  assign padl_bits_zero_124 = 0;
  assign padl_120 = { padl_bits_zero_124, padl_bits_121 };
  wire [92-1:0] padl_125;
  wire [46-1:0] padl_bits_126;
  wire [46-1:0] padl_127;
  wire [43-1:0] padl_bits_128;
  wire [43-1:0] param_129;
  assign param_129 = p_to_tau;
  assign padl_bits_128 = param_129;
  wire [3-1:0] padl_bits_zero_130;
  assign padl_bits_zero_130 = 0;
  assign padl_127 = { padl_bits_zero_130, padl_bits_128 };
  assign padl_bits_126 = padl_127;
  wire [46-1:0] padl_bits_zero_131;
  assign padl_bits_zero_131 = 0;
  assign padl_125 = { padl_bits_zero_131, padl_bits_126 };
  assign truncval_119 = padl_120 * padl_125;
  assign truncR_118 = truncval_119[85:0];
  assign toSInt_imm_117 = { toSInt_116, truncR_118[85:34] };
  assign padl_bits_115 = toSInt_imm_117;
  assign padl_114 = { { 1{ padl_bits_115[52] } }, padl_bits_115 };
  wire [54-1:0] padr_132;
  wire [11-1:0] padr_bits_133;
  assign padr_bits_133 = 0;
  wire [43-1:0] padl_134;
  wire [42-1:0] padl_bits_135;
  wire [1-1:0] toSInt_136;
  assign toSInt_136 = 0;
  wire [42-1:0] toSInt_imm_137;
  wire [41-1:0] param_138;
  assign param_138 = const_tau;
  assign toSInt_imm_137 = { toSInt_136, param_138 };
  assign padl_bits_135 = toSInt_imm_137;
  assign padl_134 = { { 1{ padl_bits_135[41] } }, padl_bits_135 };
  assign padr_132 = { padl_134, padr_bits_133 };
  assign toUsInt_95 = padr_96 + padl_114 + padr_132;
  assign truncval_94 = toUsInt_95[50:0];
  assign truncR_93 = truncval_94[51:0];
  assign tau = truncR_93[51:1];
  wire [13-1:0] truncR_139;
  wire [14-1:0] truncval_140;
  wire [15-1:0] toUsInt_141;
  wire [35-1:0] truncR_142;
  assign truncR_142 = o;
  wire [15-1:0] truncR_shift_143;
  assign truncR_shift_143 = truncR_142 >>> 20;
  wire [15-1:0] truncR_imm_144;
  assign truncR_imm_144 = (truncR_142[34])? truncR_shift_143[14:0] : truncR_142[34:20];
  assign toUsInt_141 = truncR_imm_144;
  assign truncval_140 = toUsInt_141[11:0];
  assign truncR_139 = truncval_140[12:0];
  wire [36-1:0] padl_145;
  wire [13-1:0] padl_bits_146;
  wire [36-1:0] truncR_147;
  wire [72-1:0] truncR_148;
  wire [105-1:0] truncval_149;
  wire [105-1:0] padl_150;
  wire [52-1:0] padl_bits_151;
  wire [52-1:0] padl_152;
  wire [23-1:0] padl_bits_153;
  wire [23-1:0] neg_imm_154;
  wire [23-1:0] padr_155;
  wire [8-1:0] padr_bits_156;
  assign padr_bits_156 = 0;
  wire [35-1:0] truncR_157;
  assign truncR_157 = o;
  wire [15-1:0] truncR_shift_158;
  assign truncR_shift_158 = truncR_157 >>> 20;
  wire [15-1:0] truncR_imm_159;
  assign truncR_imm_159 = (truncR_157[34])? truncR_shift_158[14:0] : truncR_157[34:20];
  assign padr_155 = { truncR_imm_159, padr_bits_156 };
  assign neg_imm_154 = -padr_155;
  assign padl_bits_153 = neg_imm_154;
  assign padl_152 = { { 29{ padl_bits_153[22] } }, padl_bits_153 };
  assign padl_bits_151 = padl_152;
  assign padl_150 = { { 53{ padl_bits_151[51] } }, padl_bits_151 };
  wire [105-1:0] padl_160;
  wire [52-1:0] padl_bits_161;
  wire [52-1:0] padr_162;
  wire [18-1:0] padr_bits_163;
  assign padr_bits_163 = 0;
  wire [1-1:0] toSInt_164;
  assign toSInt_164 = 0;
  wire [34-1:0] toSInt_imm_165;
  wire [51-1:0] truncval_166;
  assign truncval_166 = 52'd2251799813685248 / tau;
  assign toSInt_imm_165 = { toSInt_164, truncval_166[32:0] };
  assign padr_162 = { toSInt_imm_165, padr_bits_163 };
  assign padl_bits_161 = padr_162;
  assign padl_160 = { { 53{ padl_bits_161[51] } }, padl_bits_161 };
  assign truncval_149 = padl_150 * padl_160;
  wire [72-1:0] truncval_imm_167;
  assign truncval_imm_167 = { truncval_149[104], truncval_149[70:0] };
  assign truncR_148 = truncval_imm_167;
  wire [36-1:0] truncR_shift_168;
  assign truncR_shift_168 = truncR_148 >>> 36;
  wire [36-1:0] truncR_imm_169;
  assign truncR_imm_169 = (truncR_148[71])? truncR_shift_168[35:0] : truncR_148[71:36];
  assign truncR_147 = truncR_imm_169;
  wire [13-1:0] truncR_shift_170;
  assign truncR_shift_170 = truncR_147 >>> 23;
  wire [13-1:0] truncR_imm_171;
  assign truncR_imm_171 = (truncR_147[35])? truncR_shift_170[12:0] : truncR_147[35:23];
  assign padl_bits_146 = truncR_imm_171;
  assign padl_145 = { { 23{ padl_bits_146[12] } }, padl_bits_146 };
  assign dvdt = padl_145;
  wire [35-1:0] padr_172;
  wire [20-1:0] padr_bits_173;
  assign padr_bits_173 = 0;
  wire [25-1:0] truncR_174;
  wire [25-1:0] padl_175;
  wire [23-1:0] padl_bits_176;
  wire [126-1:0] truncR_177;
  wire [196-1:0] truncval_178;
  wire [196-1:0] padl_179;
  wire [109-1:0] padl_bits_180;
  wire [109-1:0] padl_181;
  wire [74-1:0] padl_bits_182;
  wire [1-1:0] toSInt_183;
  assign toSInt_183 = 0;
  wire [74-1:0] toSInt_imm_184;
  wire [73-1:0] const_185;
  assign const_185 = 73'd944473296573;
  assign toSInt_imm_184 = { toSInt_183, const_185 };
  assign padl_bits_182 = toSInt_imm_184;
  assign padl_181 = { { 35{ padl_bits_182[73] } }, padl_bits_182 };
  assign padl_bits_180 = padl_181;
  assign padl_179 = { { 87{ padl_bits_180[108] } }, padl_bits_180 };
  wire [196-1:0] padl_186;
  wire [109-1:0] padl_bits_187;
  wire [109-1:0] padr_188;
  wire [73-1:0] padr_bits_189;
  assign padr_bits_189 = 0;
  assign padr_188 = { dvdt, padr_bits_189 };
  assign padl_bits_187 = padr_188;
  assign padl_186 = { { 87{ padl_bits_187[108] } }, padl_bits_187 };
  assign truncval_178 = padl_179 * padl_186;
  wire [126-1:0] truncval_imm_190;
  assign truncval_imm_190 = { truncval_178[195], truncval_178[124:0] };
  assign truncR_177 = truncval_imm_190;
  wire [23-1:0] truncR_shift_191;
  assign truncR_shift_191 = truncR_177 >>> 103;
  wire [23-1:0] truncR_imm_192;
  assign truncR_imm_192 = (truncR_177[125])? truncR_shift_191[22:0] : truncR_177[125:103];
  assign padl_bits_176 = truncR_imm_192;
  assign padl_175 = { { 2{ padl_bits_176[22] } }, padl_bits_176 };
  assign truncR_174 = padl_175;
  wire [15-1:0] truncR_shift_193;
  assign truncR_shift_193 = truncR_174 >>> 10;
  wire [15-1:0] truncR_imm_194;
  assign truncR_imm_194 = (truncR_174[24])? truncR_shift_193[14:0] : truncR_174[24:10];
  assign padr_172 = { truncR_imm_194, padr_bits_173 };
  wire [32-1:0] padl_195;
  wire [2-1:0] padl_bits_196;
  wire [13-1:0] truncR_197;
  wire [23-1:0] truncR_198;
  wire [114-1:0] truncR_199;
  wire [182-1:0] truncval_200;
  wire [182-1:0] padl_201;
  wire [91-1:0] padl_bits_202;
  wire [91-1:0] padl_203;
  wire [58-1:0] padl_bits_204;
  wire [98-1:0] truncR_205;
  wire [105-1:0] truncval_206;
  wire [105-1:0] padl_207;
  wire [52-1:0] padl_bits_208;
  wire [52-1:0] padr_209;
  wire [41-1:0] padr_bits_210;
  assign padr_bits_210 = 0;
  wire [1-1:0] toSInt_211;
  assign toSInt_211 = 0;
  wire [11-1:0] toSInt_imm_212;
  assign toSInt_imm_212 = { toSInt_211, n };
  assign padr_209 = { toSInt_imm_212, padr_bits_210 };
  assign padl_bits_208 = padr_209;
  assign padl_207 = { { 53{ padl_bits_208[51] } }, padl_bits_208 };
  wire [105-1:0] padl_213;
  wire [52-1:0] padl_bits_214;
  wire [52-1:0] padl_215;
  wire [50-1:0] padl_bits_216;
  wire [50-1:0] param_217;
  assign param_217 = n_to_response_time_lh;
  assign padl_bits_216 = param_217;
  assign padl_215 = { { 2{ padl_bits_216[49] } }, padl_bits_216 };
  assign padl_bits_214 = padl_215;
  assign padl_213 = { { 53{ padl_bits_214[51] } }, padl_bits_214 };
  assign truncval_206 = padl_207 * padl_213;
  wire [98-1:0] truncval_imm_218;
  assign truncval_imm_218 = { truncval_206[104], truncval_206[96:0] };
  assign truncR_205 = truncval_imm_218;
  wire [58-1:0] truncR_shift_219;
  assign truncR_shift_219 = truncR_205 >>> 40;
  wire [58-1:0] truncR_imm_220;
  assign truncR_imm_220 = (truncR_205[97])? truncR_shift_219[57:0] : truncR_205[97:40];
  wire [58-1:0] padr_221;
  wire [1-1:0] padr_bits_222;
  assign padr_bits_222 = 0;
  wire [94-1:0] truncR_223;
  wire [101-1:0] truncval_224;
  wire [101-1:0] padl_225;
  wire [50-1:0] padl_bits_226;
  wire [50-1:0] padr_227;
  wire [39-1:0] padr_bits_228;
  assign padr_bits_228 = 0;
  wire [1-1:0] toSInt_229;
  assign toSInt_229 = 0;
  wire [11-1:0] toSInt_imm_230;
  assign toSInt_imm_230 = { toSInt_229, p };
  assign padr_227 = { toSInt_imm_230, padr_bits_228 };
  assign padl_bits_226 = padr_227;
  assign padl_225 = { { 51{ padl_bits_226[49] } }, padl_bits_226 };
  wire [101-1:0] padl_231;
  wire [50-1:0] padl_bits_232;
  wire [50-1:0] padl_233;
  wire [48-1:0] padl_bits_234;
  wire [48-1:0] param_235;
  assign param_235 = p_to_response_time_lh;
  assign padl_bits_234 = param_235;
  assign padl_233 = { { 2{ padl_bits_234[47] } }, padl_bits_234 };
  assign padl_bits_232 = padl_233;
  assign padl_231 = { { 51{ padl_bits_232[49] } }, padl_bits_232 };
  assign truncval_224 = padl_225 * padl_231;
  wire [94-1:0] truncval_imm_236;
  assign truncval_imm_236 = { truncval_224[100], truncval_224[92:0] };
  assign truncR_223 = truncval_imm_236;
  wire [57-1:0] truncR_shift_237;
  assign truncR_shift_237 = truncR_223 >>> 37;
  wire [57-1:0] truncR_imm_238;
  assign truncR_imm_238 = (truncR_223[93])? truncR_shift_237[56:0] : truncR_223[93:37];
  assign padr_221 = { truncR_imm_238, padr_bits_222 };
  wire [58-1:0] padr_239;
  wire [13-1:0] padr_bits_240;
  assign padr_bits_240 = 0;
  wire [45-1:0] padl_241;
  wire [44-1:0] padl_bits_242;
  wire [1-1:0] toSInt_243;
  assign toSInt_243 = 0;
  wire [44-1:0] toSInt_imm_244;
  wire [43-1:0] param_245;
  assign param_245 = const_response_time_lh;
  assign toSInt_imm_244 = { toSInt_243, param_245 };
  assign padl_bits_242 = toSInt_imm_244;
  assign padl_241 = { { 1{ padl_bits_242[43] } }, padl_bits_242 };
  assign padr_239 = { padl_241, padr_bits_240 };
  assign padl_bits_204 = truncR_imm_220 + padr_221 + padr_239;
  assign padl_203 = { { 33{ padl_bits_204[57] } }, padl_bits_204 };
  assign padl_bits_202 = padl_203;
  assign padl_201 = { { 91{ padl_bits_202[90] } }, padl_bits_202 };
  wire [182-1:0] padl_246;
  wire [91-1:0] padl_bits_247;
  wire [91-1:0] padr_248;
  wire [50-1:0] padr_bits_249;
  assign padr_bits_249 = 0;
  wire [1-1:0] toSInt_250;
  assign toSInt_250 = 0;
  wire [41-1:0] toSInt_imm_251;
  wire [40-1:0] const_252;
  assign const_252 = 40'd640000000000;
  assign toSInt_imm_251 = { toSInt_250, const_252 };
  assign padr_248 = { toSInt_imm_251, padr_bits_249 };
  assign padl_bits_247 = padr_248;
  assign padl_246 = { { 91{ padl_bits_247[90] } }, padl_bits_247 };
  assign truncval_200 = padl_201 * padl_246;
  assign truncR_199 = truncval_200[113:0];
  assign truncR_198 = truncR_199[113:91];
  assign truncR_197 = truncR_198[22:10];
  assign padl_bits_196 = truncR_197[12:11];
  wire [30-1:0] padl_bits_zero_253;
  assign padl_bits_zero_253 = 0;
  assign padl_195 = { padl_bits_zero_253, padl_bits_196 };
  assign wait_time_lh = padl_195;
  wire [35-1:0] padr_254;
  wire [20-1:0] padr_bits_255;
  assign padr_bits_255 = 0;
  wire [54-1:0] truncR_256;
  wire [54-1:0] padl_257;
  wire [50-1:0] padl_bits_258;
  wire [1-1:0] toSInt_259;
  assign toSInt_259 = 0;
  wire [50-1:0] toSInt_imm_260;
  wire [49-1:0] const_261;
  assign const_261 = 49'd562949953421;
  assign toSInt_imm_260 = { toSInt_259, const_261 };
  assign padl_bits_258 = toSInt_imm_260;
  assign padl_257 = { { 4{ padl_bits_258[49] } }, padl_bits_258 };
  assign truncR_256 = padl_257;
  wire [15-1:0] truncR_shift_262;
  assign truncR_shift_262 = truncR_256 >>> 39;
  wire [15-1:0] truncR_imm_263;
  assign truncR_imm_263 = (truncR_256[53])? truncR_shift_262[14:0] : truncR_256[53:39];
  assign padr_254 = { truncR_imm_263, padr_bits_255 };
  wire [13-1:0] truncR_264;
  wire [14-1:0] truncval_265;
  wire [15-1:0] toUsInt_266;
  wire [35-1:0] truncR_267;
  assign truncR_267 = o;
  wire [15-1:0] truncR_shift_268;
  assign truncR_shift_268 = truncR_267 >>> 20;
  wire [15-1:0] truncR_imm_269;
  assign truncR_imm_269 = (truncR_267[34])? truncR_shift_268[14:0] : truncR_267[34:20];
  assign toUsInt_266 = truncR_imm_269;
  assign truncval_265 = toUsInt_266[11:0];
  assign truncR_264 = truncval_265[12:0];
  wire [59-1:0] padr_270;
  wire [3-1:0] padr_bits_271;
  assign padr_bits_271 = 0;
  wire [57-1:0] truncval_272;
  wire [58-1:0] toUsInt_273;
  wire [58-1:0] padr_274;
  wire [3-1:0] padr_bits_275;
  assign padr_bits_275 = 0;
  wire [55-1:0] padl_276;
  wire [54-1:0] padl_bits_277;
  wire [1-1:0] toSInt_278;
  assign toSInt_278 = 0;
  wire [54-1:0] toSInt_imm_279;
  wire [88-1:0] truncR_280;
  wire [94-1:0] truncval_281;
  wire [94-1:0] padl_282;
  wire [47-1:0] padl_bits_283;
  wire [47-1:0] padr_284;
  wire [37-1:0] padr_bits_285;
  assign padr_bits_285 = 0;
  assign padr_284 = { n, padr_bits_285 };
  assign padl_bits_283 = padr_284;
  wire [47-1:0] padl_bits_zero_286;
  assign padl_bits_zero_286 = 0;
  assign padl_282 = { padl_bits_zero_286, padl_bits_283 };
  wire [94-1:0] padl_287;
  wire [47-1:0] padl_bits_288;
  wire [47-1:0] padl_289;
  wire [44-1:0] padl_bits_290;
  wire [44-1:0] param_291;
  assign param_291 = n_to_tau_lh;
  assign padl_bits_290 = param_291;
  wire [3-1:0] padl_bits_zero_292;
  assign padl_bits_zero_292 = 0;
  assign padl_289 = { padl_bits_zero_292, padl_bits_290 };
  assign padl_bits_288 = padl_289;
  wire [47-1:0] padl_bits_zero_293;
  assign padl_bits_zero_293 = 0;
  assign padl_287 = { padl_bits_zero_293, padl_bits_288 };
  assign truncval_281 = padl_282 * padl_287;
  assign truncR_280 = truncval_281[87:0];
  assign toSInt_imm_279 = { toSInt_278, truncR_280[87:35] };
  assign padl_bits_277 = toSInt_imm_279;
  assign padl_276 = { { 1{ padl_bits_277[53] } }, padl_bits_277 };
  assign padr_274 = { padl_276, padr_bits_275 };
  wire [96-1:0] truncR_294;
  wire [103-1:0] truncval_295;
  wire [103-1:0] padl_296;
  wire [51-1:0] padl_bits_297;
  wire [51-1:0] padr_298;
  wire [40-1:0] padr_bits_299;
  assign padr_bits_299 = 0;
  wire [1-1:0] toSInt_300;
  assign toSInt_300 = 0;
  wire [11-1:0] toSInt_imm_301;
  assign toSInt_imm_301 = { toSInt_300, p };
  assign padr_298 = { toSInt_imm_301, padr_bits_299 };
  assign padl_bits_297 = padr_298;
  assign padl_296 = { { 52{ padl_bits_297[50] } }, padl_bits_297 };
  wire [103-1:0] padl_302;
  wire [51-1:0] padl_bits_303;
  wire [51-1:0] padl_304;
  wire [49-1:0] padl_bits_305;
  wire [49-1:0] param_306;
  assign param_306 = p_to_tau_lh;
  assign padl_bits_305 = param_306;
  assign padl_304 = { { 2{ padl_bits_305[48] } }, padl_bits_305 };
  assign padl_bits_303 = padl_304;
  assign padl_302 = { { 52{ padl_bits_303[50] } }, padl_bits_303 };
  assign truncval_295 = padl_296 * padl_302;
  wire [96-1:0] truncval_imm_307;
  assign truncval_imm_307 = { truncval_295[102], truncval_295[94:0] };
  assign truncR_294 = truncval_imm_307;
  wire [58-1:0] truncR_shift_308;
  assign truncR_shift_308 = truncR_294 >>> 38;
  wire [58-1:0] truncR_imm_309;
  assign truncR_imm_309 = (truncR_294[95])? truncR_shift_308[57:0] : truncR_294[95:38];
  wire [58-1:0] padr_310;
  wire [13-1:0] padr_bits_311;
  assign padr_bits_311 = 0;
  wire [45-1:0] padl_312;
  wire [44-1:0] padl_bits_313;
  wire [1-1:0] toSInt_314;
  assign toSInt_314 = 0;
  wire [44-1:0] toSInt_imm_315;
  wire [43-1:0] param_316;
  assign param_316 = const_tau_lh;
  assign toSInt_imm_315 = { toSInt_314, param_316 };
  assign padl_bits_313 = toSInt_imm_315;
  assign padl_312 = { { 1{ padl_bits_313[43] } }, padl_bits_313 };
  assign padr_310 = { padl_312, padr_bits_311 };
  assign toUsInt_273 = padr_274 + truncR_imm_309 + padr_310;
  assign truncval_272 = toUsInt_273[54:0];
  assign padr_270 = { truncval_272[55:0], padr_bits_271 };
  assign tau_lh = padr_270;
  wire [33-1:0] truncR_317;
  wire [34-1:0] truncval_318;
  wire [35-1:0] toUsInt_319;
  assign toUsInt_319 = o;
  assign truncval_318 = toUsInt_319[31:0];
  assign truncR_317 = truncval_318[32:0];
  wire [37-1:0] padl_320;
  wire [13-1:0] padl_bits_321;
  wire [37-1:0] truncR_322;
  wire [113-1:0] truncR_323;
  wire [145-1:0] truncval_324;
  wire [145-1:0] padl_325;
  wire [72-1:0] padl_bits_326;
  wire [72-1:0] padl_327;
  wire [43-1:0] padl_bits_328;
  wire [43-1:0] padl_329;
  wire [41-1:0] padl_bits_330;
  wire [1-1:0] toSInt_331;
  assign toSInt_331 = 0;
  wire [41-1:0] toSInt_imm_332;
  wire [40-1:0] const_333;
  assign const_333 = 40'd907097092915;
  assign toSInt_imm_332 = { toSInt_331, const_333 };
  assign padl_bits_330 = toSInt_imm_332;
  assign padl_329 = { { 2{ padl_bits_330[40] } }, padl_bits_330 };
  wire [43-1:0] padr_334;
  wire [8-1:0] padr_bits_335;
  assign padr_bits_335 = 0;
  assign padr_334 = { o, padr_bits_335 };
  assign padl_bits_328 = padl_329 - padr_334;
  assign padl_327 = { { 29{ padl_bits_328[42] } }, padl_bits_328 };
  assign padl_bits_326 = padl_327;
  assign padl_325 = { { 73{ padl_bits_326[71] } }, padl_bits_326 };
  wire [145-1:0] padl_336;
  wire [72-1:0] padl_bits_337;
  wire [72-1:0] padr_338;
  wire [38-1:0] padr_bits_339;
  assign padr_bits_339 = 0;
  wire [1-1:0] toSInt_340;
  assign toSInt_340 = 0;
  wire [34-1:0] toSInt_imm_341;
  wire [59-1:0] truncval_342;
  assign truncval_342 = 60'd576460752303423488 / tau_lh;
  assign toSInt_imm_341 = { toSInt_340, truncval_342[32:0] };
  assign padr_338 = { toSInt_imm_341, padr_bits_339 };
  assign padl_bits_337 = padr_338;
  assign padl_336 = { { 73{ padl_bits_337[71] } }, padl_bits_337 };
  assign truncval_324 = padl_325 * padl_336;
  wire [113-1:0] truncval_imm_343;
  assign truncval_imm_343 = { truncval_324[144], truncval_324[111:0] };
  assign truncR_323 = truncval_imm_343;
  wire [37-1:0] truncR_shift_344;
  assign truncR_shift_344 = truncR_323 >>> 76;
  wire [37-1:0] truncR_imm_345;
  assign truncR_imm_345 = (truncR_323[112])? truncR_shift_344[36:0] : truncR_323[112:76];
  assign truncR_322 = truncR_imm_345;
  wire [13-1:0] truncR_shift_346;
  assign truncR_shift_346 = truncR_322 >>> 24;
  wire [13-1:0] truncR_imm_347;
  assign truncR_imm_347 = (truncR_322[36])? truncR_shift_346[12:0] : truncR_322[36:24];
  assign padl_bits_321 = truncR_imm_347;
  assign padl_320 = { { 24{ padl_bits_321[12] } }, padl_bits_321 };
  assign dodt = padl_320;
  wire [35-1:0] padr_348;
  wire [10-1:0] padr_bits_349;
  assign padr_bits_349 = 0;
  wire [25-1:0] padl_350;
  wire [23-1:0] padl_bits_351;
  wire [125-1:0] truncR_352;
  wire [197-1:0] truncval_353;
  wire [197-1:0] padl_354;
  wire [110-1:0] padl_bits_355;
  wire [110-1:0] padl_356;
  wire [74-1:0] padl_bits_357;
  wire [1-1:0] toSInt_358;
  assign toSInt_358 = 0;
  wire [74-1:0] toSInt_imm_359;
  wire [73-1:0] const_360;
  assign const_360 = 73'd944473296573;
  assign toSInt_imm_359 = { toSInt_358, const_360 };
  assign padl_bits_357 = toSInt_imm_359;
  assign padl_356 = { { 36{ padl_bits_357[73] } }, padl_bits_357 };
  assign padl_bits_355 = padl_356;
  assign padl_354 = { { 87{ padl_bits_355[109] } }, padl_bits_355 };
  wire [197-1:0] padl_361;
  wire [110-1:0] padl_bits_362;
  wire [110-1:0] padr_363;
  wire [73-1:0] padr_bits_364;
  assign padr_bits_364 = 0;
  assign padr_363 = { dodt, padr_bits_364 };
  assign padl_bits_362 = padr_363;
  assign padl_361 = { { 87{ padl_bits_362[109] } }, padl_bits_362 };
  assign truncval_353 = padl_354 * padl_361;
  wire [125-1:0] truncval_imm_365;
  assign truncval_imm_365 = { truncval_353[196], truncval_353[123:0] };
  assign truncR_352 = truncval_imm_365;
  wire [23-1:0] truncR_shift_366;
  assign truncR_shift_366 = truncR_352 >>> 102;
  wire [23-1:0] truncR_imm_367;
  assign truncR_imm_367 = (truncR_352[124])? truncR_shift_366[22:0] : truncR_352[124:102];
  assign padl_bits_351 = truncR_imm_367;
  assign padl_350 = { { 2{ padl_bits_351[22] } }, padl_bits_351 };
  assign padr_348 = { padl_350, padr_bits_349 };
  assign out = (fsm == 0)? truncR_10[12:3] : truncR_87[12:3];

  always @(posedge clk) begin
    prev_sys_clk <= sys_clk;
  end

  localparam fsm_1 = 1;
  localparam fsm_2 = 2;
  localparam fsm_3 = 3;
  localparam fsm_4 = 4;

  always @(posedge clk) begin
    if(reset) begin
      fsm <= fsm_init;
    end else begin
      case(fsm)
        fsm_init: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_0;
          end
          if(~prev_sys_clk & sys_clk & ((n > p) & (n <= 10'd512))) begin
            fsm <= fsm_1;
          end 
        end
        fsm_1: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_77;
          end
          if(state_cycle_counter > wait_time) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time) begin
            fsm <= fsm_2;
          end 
        end
        fsm_2: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= o + padr_172;
          end
          if(prev_sys_clk & ~sys_clk) begin
            fsm <= fsm_3;
          end 
        end
        fsm_3: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_254;
          end
          if(state_cycle_counter > wait_time_lh) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time_lh) begin
            fsm <= fsm_4;
          end 
        end
        fsm_4: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= o + padr_348;
          end
          if((o > 35'd3532610600) & (o <= 35'd17179869184)) begin
            fsm <= fsm_init;
          end 
        end
      endcase
    end
  end


endmodule


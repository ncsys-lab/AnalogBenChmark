

module voltage_controlled_oscillator #
(
  parameter gain = 1024,
  parameter rest_frec = 1638
)
(
  input clk,
  input reset,
  input [10-1:0] input_voltage_real,
  output [31-1:0] output_clock_real
);

  reg [31-1:0] x;
  reg [31-1:0] v;
  reg [10-1:0] input_voltage_prev;
  wire [26-1:0] dwdt;
  wire [26-1:0] dvdt;
  wire [26-1:0] dxdt;
  reg [10-1:0] prev_input_voltage_real;
  wire [83-1:0] truncR_0;
  wire [95-1:0] truncval_1;
  wire [95-1:0] padl_2;
  wire [47-1:0] padl_bits_3;
  wire [47-1:0] padr_4;
  wire [25-1:0] padr_bits_5;
  assign padr_bits_5 = 0;
  wire [22-1:0] padl_6;
  wire [10-1:0] padl_bits_7;
  assign padl_bits_7 = input_voltage_real - input_voltage_prev;
  wire [12-1:0] padl_bits_zero_8;
  assign padl_bits_zero_8 = 0;
  assign padl_6 = { padl_bits_zero_8, padl_bits_7 };
  assign padr_4 = { padl_6, padr_bits_5 };
  assign padl_bits_3 = padr_4;
  wire [48-1:0] padl_bits_zero_9;
  assign padl_bits_zero_9 = 0;
  assign padl_2 = { padl_bits_zero_9, padl_bits_3 };
  wire [95-1:0] padl_10;
  wire [47-1:0] padl_bits_11;
  wire [47-1:0] const_12;
  assign const_12 = 47'd85899345920000;
  assign padl_bits_11 = const_12;
  wire [48-1:0] padl_bits_zero_13;
  assign padl_bits_zero_13 = 0;
  assign padl_10 = { padl_bits_zero_13, padl_bits_11 };
  assign truncval_1 = padl_2 * padl_10;
  wire [83-1:0] truncval_imm_14;
  assign truncval_imm_14 = { truncval_1[94], truncval_1[81:0] };
  assign truncR_0 = truncval_imm_14;
  wire [26-1:0] truncR_shift_15;
  assign truncR_shift_15 = truncR_0 >>> 57;
  wire [26-1:0] truncR_imm_16;
  assign truncR_imm_16 = (truncR_0[82])? truncR_shift_15[25:0] : truncR_0[82:57];
  assign dwdt = truncR_imm_16;
  wire [31-1:0] truncR_17;
  wire [31-1:0] padl_18;
  wire [26-1:0] padl_bits_19;
  wire [57-1:0] truncR_20;
  wire [63-1:0] truncval_21;
  wire [63-1:0] padl_22;
  wire [31-1:0] padl_bits_23;
  wire [31-1:0] padr_24;
  wire [4-1:0] padr_bits_25;
  assign padr_bits_25 = 0;
  wire [27-1:0] padl_26;
  wire [26-1:0] padl_bits_27;
  wire [26-1:0] neg_imm_28;
  wire [46-1:0] truncR_29;
  wire [53-1:0] truncval_30;
  wire [53-1:0] padl_31;
  wire [26-1:0] padl_bits_32;
  wire [50-1:0] truncR_33;
  wire [51-1:0] truncval_34;
  wire [51-1:0] padl_35;
  wire [25-1:0] padl_bits_36;
  wire [25-1:0] padr_37;
  wire [2-1:0] padr_bits_38;
  assign padr_bits_38 = 0;
  wire [26-1:0] truncval_39;
  wire [26-1:0] padl_40;
  wire [13-1:0] padl_bits_41;
  wire [13-1:0] padl_42;
  wire [11-1:0] padl_bits_43;
  wire [11-1:0] param_44;
  assign param_44 = gain;
  assign padl_bits_43 = param_44;
  wire [2-1:0] padl_bits_zero_45;
  assign padl_bits_zero_45 = 0;
  assign padl_42 = { padl_bits_zero_45, padl_bits_43 };
  assign padl_bits_41 = padl_42;
  wire [13-1:0] padl_bits_zero_46;
  assign padl_bits_zero_46 = 0;
  assign padl_40 = { padl_bits_zero_46, padl_bits_41 };
  wire [26-1:0] padl_47;
  wire [13-1:0] padl_bits_48;
  wire [13-1:0] padr_49;
  wire [3-1:0] padr_bits_50;
  assign padr_bits_50 = 0;
  assign padr_49 = { input_voltage_real, padr_bits_50 };
  assign padl_bits_48 = padr_49;
  wire [13-1:0] padl_bits_zero_51;
  assign padl_bits_zero_51 = 0;
  assign padl_47 = { padl_bits_zero_51, padl_bits_48 };
  assign truncval_39 = padl_40 * padl_47;
  assign padr_37 = { truncval_39[22:0], padr_bits_38 };
  assign padl_bits_36 = padr_37;
  wire [26-1:0] padl_bits_zero_52;
  assign padl_bits_zero_52 = 0;
  assign padl_35 = { padl_bits_zero_52, padl_bits_36 };
  wire [51-1:0] padl_53;
  wire [25-1:0] padl_bits_54;
  wire [25-1:0] padr_55;
  wire [15-1:0] padr_bits_56;
  assign padr_bits_56 = 0;
  assign padr_55 = { input_voltage_real, padr_bits_56 };
  assign padl_bits_54 = padr_55;
  wire [26-1:0] padl_bits_zero_57;
  assign padl_bits_zero_57 = 0;
  assign padl_53 = { padl_bits_zero_57, padl_bits_54 };
  assign truncval_34 = padl_35 * padl_53;
  wire [50-1:0] truncval_imm_58;
  assign truncval_imm_58 = { truncval_34[50], truncval_34[48:0] };
  assign truncR_33 = truncval_imm_58;
  wire [26-1:0] truncR_shift_59;
  assign truncR_shift_59 = truncR_33 >>> 24;
  wire [26-1:0] truncR_imm_60;
  assign truncR_imm_60 = (truncR_33[49])? truncR_shift_59[25:0] : truncR_33[49:24];
  assign padl_bits_32 = truncR_imm_60;
  assign padl_31 = { { 27{ padl_bits_32[25] } }, padl_bits_32 };
  wire [53-1:0] padl_61;
  wire [26-1:0] padl_bits_62;
  wire [26-1:0] padr_63;
  wire [10-1:0] padr_bits_64;
  assign padr_bits_64 = 0;
  wire [16-1:0] padl_65;
  wire [12-1:0] padl_bits_66;
  wire [1-1:0] toSInt_67;
  assign toSInt_67 = 0;
  wire [12-1:0] toSInt_imm_68;
  wire [11-1:0] param_69;
  assign param_69 = gain;
  assign toSInt_imm_68 = { toSInt_67, param_69 };
  assign padl_bits_66 = toSInt_imm_68;
  assign padl_65 = { { 4{ padl_bits_66[11] } }, padl_bits_66 };
  assign padr_63 = { padl_65, padr_bits_64 };
  assign padl_bits_62 = padr_63;
  assign padl_61 = { { 27{ padl_bits_62[25] } }, padl_bits_62 };
  assign truncval_30 = padl_31 * padl_61;
  wire [46-1:0] truncval_imm_70;
  assign truncval_imm_70 = { truncval_30[52], truncval_30[44:0] };
  assign truncR_29 = truncval_imm_70;
  wire [26-1:0] truncR_shift_71;
  assign truncR_shift_71 = truncR_29 >>> 20;
  wire [26-1:0] truncR_imm_72;
  assign truncR_imm_72 = (truncR_29[45])? truncR_shift_71[25:0] : truncR_29[45:20];
  wire [26-1:0] padr_73;
  wire [6-1:0] padr_bits_74;
  assign padr_bits_74 = 0;
  wire [20-1:0] padl_75;
  wire [15-1:0] padl_bits_76;
  wire [1-1:0] toSInt_77;
  assign toSInt_77 = 0;
  wire [15-1:0] toSInt_imm_78;
  wire [14-1:0] param_79;
  assign param_79 = rest_frec;
  assign toSInt_imm_78 = { toSInt_77, param_79 };
  assign padl_bits_76 = toSInt_imm_78;
  assign padl_75 = { { 5{ padl_bits_76[14] } }, padl_bits_76 };
  assign padr_73 = { padl_75, padr_bits_74 };
  assign neg_imm_28 = -(truncR_imm_72 + padr_73);
  assign padl_bits_27 = neg_imm_28;
  assign padl_26 = { { 1{ padl_bits_27[25] } }, padl_bits_27 };
  assign padr_24 = { padl_26, padr_bits_25 };
  assign padl_bits_23 = padr_24;
  assign padl_22 = { { 32{ padl_bits_23[30] } }, padl_bits_23 };
  wire [63-1:0] padl_80;
  wire [31-1:0] padl_bits_81;
  assign padl_bits_81 = x;
  assign padl_80 = { { 32{ padl_bits_81[30] } }, padl_bits_81 };
  assign truncval_21 = padl_22 * padl_80;
  wire [57-1:0] truncval_imm_82;
  assign truncval_imm_82 = { truncval_21[62], truncval_21[55:0] };
  assign truncR_20 = truncval_imm_82;
  wire [26-1:0] truncR_shift_83;
  assign truncR_shift_83 = truncR_20 >>> 31;
  wire [26-1:0] truncR_imm_84;
  assign truncR_imm_84 = (truncR_20[56])? truncR_shift_83[25:0] : truncR_20[56:31];
  assign padl_bits_19 = truncR_imm_84;
  assign padl_18 = { { 5{ padl_bits_19[25] } }, padl_bits_19 };
  wire [31-1:0] padr_85;
  wire [5-1:0] padr_bits_86;
  assign padr_bits_86 = 0;
  wire [62-1:0] truncR_87;
  wire [83-1:0] truncval_88;
  wire [83-1:0] padl_89;
  wire [41-1:0] padl_bits_90;
  wire [41-1:0] padr_91;
  wire [15-1:0] padr_bits_92;
  assign padr_bits_92 = 0;
  wire [67-1:0] truncR_93;
  wire [89-1:0] truncval_94;
  wire [89-1:0] padl_95;
  wire [44-1:0] padl_bits_96;
  wire [44-1:0] padl_97;
  wire [26-1:0] padl_bits_98;
  wire [1-1:0] toSInt_99;
  assign toSInt_99 = 0;
  wire [26-1:0] toSInt_imm_100;
  wire [50-1:0] truncR_101;
  wire [52-1:0] truncval_102;
  wire [52-1:0] padl_103;
  wire [26-1:0] padl_bits_104;
  wire [26-1:0] padl_105;
  wire [25-1:0] padl_bits_106;
  wire [25-1:0] padr_107;
  wire [22-1:0] padr_bits_108;
  assign padr_bits_108 = 0;
  wire [49-1:0] truncval_109;
  wire [49-1:0] padr_110;
  wire [24-1:0] padr_bits_111;
  assign padr_bits_111 = 0;
  wire [25-1:0] padr_112;
  wire [2-1:0] padr_bits_113;
  assign padr_bits_113 = 0;
  wire [26-1:0] truncval_114;
  wire [26-1:0] padl_115;
  wire [13-1:0] padl_bits_116;
  wire [13-1:0] padl_117;
  wire [11-1:0] padl_bits_118;
  wire [11-1:0] param_119;
  assign param_119 = gain;
  assign padl_bits_118 = param_119;
  wire [2-1:0] padl_bits_zero_120;
  assign padl_bits_zero_120 = 0;
  assign padl_117 = { padl_bits_zero_120, padl_bits_118 };
  assign padl_bits_116 = padl_117;
  wire [13-1:0] padl_bits_zero_121;
  assign padl_bits_zero_121 = 0;
  assign padl_115 = { padl_bits_zero_121, padl_bits_116 };
  wire [26-1:0] padl_122;
  wire [13-1:0] padl_bits_123;
  wire [13-1:0] padr_124;
  wire [3-1:0] padr_bits_125;
  assign padr_bits_125 = 0;
  assign padr_124 = { input_voltage_real, padr_bits_125 };
  assign padl_bits_123 = padr_124;
  wire [13-1:0] padl_bits_zero_126;
  assign padl_bits_zero_126 = 0;
  assign padl_122 = { padl_bits_zero_126, padl_bits_123 };
  assign truncval_114 = padl_115 * padl_122;
  assign padr_112 = { truncval_114[22:0], padr_bits_113 };
  assign padr_110 = { padr_112, padr_bits_111 };
  wire [49-1:0] padl_127;
  wire [47-1:0] padl_bits_128;
  wire [47-1:0] const_129;
  assign const_129 = 47'd70368744177664;
  assign padl_bits_128 = const_129;
  wire [2-1:0] padl_bits_zero_130;
  assign padl_bits_zero_130 = 0;
  assign padl_127 = { padl_bits_zero_130, padl_bits_128 };
  assign truncval_109 = 50'd562949953421312 / (padr_110 + padl_127);
  assign padr_107 = { truncval_109[2:0], padr_bits_108 };
  assign padl_bits_106 = padr_107;
  wire [1-1:0] padl_bits_zero_131;
  assign padl_bits_zero_131 = 0;
  assign padl_105 = { padl_bits_zero_131, padl_bits_106 };
  assign padl_bits_104 = padl_105;
  wire [26-1:0] padl_bits_zero_132;
  assign padl_bits_zero_132 = 0;
  assign padl_103 = { padl_bits_zero_132, padl_bits_104 };
  wire [52-1:0] padl_133;
  wire [26-1:0] padl_bits_134;
  wire [26-1:0] padr_135;
  wire [15-1:0] padr_bits_136;
  assign padr_bits_136 = 0;
  wire [11-1:0] param_137;
  assign param_137 = gain;
  assign padr_135 = { param_137, padr_bits_136 };
  assign padl_bits_134 = padr_135;
  wire [26-1:0] padl_bits_zero_138;
  assign padl_bits_zero_138 = 0;
  assign padl_133 = { padl_bits_zero_138, padl_bits_134 };
  assign truncval_102 = padl_103 * padl_133;
  assign truncR_101 = truncval_102[49:0];
  assign toSInt_imm_100 = { toSInt_99, truncR_101[49:25] };
  assign padl_bits_98 = toSInt_imm_100;
  assign padl_97 = { { 18{ padl_bits_98[25] } }, padl_bits_98 };
  assign padl_bits_96 = padl_97;
  assign padl_95 = { { 45{ padl_bits_96[43] } }, padl_bits_96 };
  wire [89-1:0] padl_139;
  wire [44-1:0] padl_bits_140;
  wire [44-1:0] padr_141;
  wire [18-1:0] padr_bits_142;
  assign padr_bits_142 = 0;
  assign padr_141 = { dwdt, padr_bits_142 };
  assign padl_bits_140 = padr_141;
  assign padl_139 = { { 45{ padl_bits_140[43] } }, padl_bits_140 };
  assign truncval_94 = padl_95 * padl_139;
  wire [67-1:0] truncval_imm_143;
  assign truncval_imm_143 = { truncval_94[88], truncval_94[65:0] };
  assign truncR_93 = truncval_imm_143;
  wire [26-1:0] truncR_shift_144;
  assign truncR_shift_144 = truncR_93 >>> 41;
  wire [26-1:0] truncR_imm_145;
  assign truncR_imm_145 = (truncR_93[66])? truncR_shift_144[25:0] : truncR_93[66:41];
  assign padr_91 = { truncR_imm_145, padr_bits_92 };
  assign padl_bits_90 = padr_91;
  assign padl_89 = { { 42{ padl_bits_90[40] } }, padl_bits_90 };
  wire [83-1:0] padl_146;
  wire [41-1:0] padl_bits_147;
  wire [41-1:0] padl_148;
  wire [31-1:0] padl_bits_149;
  assign padl_bits_149 = v;
  assign padl_148 = { { 10{ padl_bits_149[30] } }, padl_bits_149 };
  assign padl_bits_147 = padl_148;
  assign padl_146 = { { 42{ padl_bits_147[40] } }, padl_bits_147 };
  assign truncval_88 = padl_89 * padl_146;
  wire [62-1:0] truncval_imm_150;
  assign truncval_imm_150 = { truncval_88[82], truncval_88[60:0] };
  assign truncR_87 = truncval_imm_150;
  wire [26-1:0] truncR_shift_151;
  assign truncR_shift_151 = truncR_87 >>> 36;
  wire [26-1:0] truncR_imm_152;
  assign truncR_imm_152 = (truncR_87[61])? truncR_shift_151[25:0] : truncR_87[61:36];
  assign padr_85 = { truncR_imm_152, padr_bits_86 };
  assign truncR_17 = padl_18 + padr_85;
  wire [26-1:0] truncR_shift_153;
  assign truncR_shift_153 = truncR_17 >>> 5;
  wire [26-1:0] truncR_imm_154;
  assign truncR_imm_154 = (truncR_17[30])? truncR_shift_153[25:0] : truncR_17[30:5];
  assign dvdt = truncR_imm_154;
  wire [31-1:0] truncR_155;
  assign truncR_155 = v;
  wire [26-1:0] truncR_shift_156;
  assign truncR_shift_156 = truncR_155 >>> 5;
  wire [26-1:0] truncR_imm_157;
  assign truncR_imm_157 = (truncR_155[30])? truncR_shift_156[25:0] : truncR_155[30:5];
  assign dxdt = truncR_imm_157;
  assign output_clock_real = x;
  wire [33-1:0] truncR_158;
  wire [33-1:0] padl_159;
  wire [28-1:0] padl_bits_160;
  wire [122-1:0] truncR_161;
  wire [149-1:0] truncval_162;
  wire [149-1:0] padl_163;
  wire [74-1:0] padl_bits_164;
  wire [74-1:0] padl_165;
  wire [61-1:0] padl_bits_166;
  wire [1-1:0] toSInt_167;
  assign toSInt_167 = 0;
  wire [61-1:0] toSInt_imm_168;
  wire [60-1:0] const_169;
  assign const_169 = 60'd57646075230342;
  assign toSInt_imm_168 = { toSInt_167, const_169 };
  assign padl_bits_166 = toSInt_imm_168;
  assign padl_165 = { { 13{ padl_bits_166[60] } }, padl_bits_166 };
  assign padl_bits_164 = padl_165;
  assign padl_163 = { { 75{ padl_bits_164[73] } }, padl_bits_164 };
  wire [149-1:0] padl_170;
  wire [74-1:0] padl_bits_171;
  wire [74-1:0] padr_172;
  wire [48-1:0] padr_bits_173;
  assign padr_bits_173 = 0;
  assign padr_172 = { dvdt, padr_bits_173 };
  assign padl_bits_171 = padr_172;
  assign padl_170 = { { 75{ padl_bits_171[73] } }, padl_bits_171 };
  assign truncval_162 = padl_163 * padl_170;
  wire [122-1:0] truncval_imm_174;
  assign truncval_imm_174 = { truncval_162[148], truncval_162[120:0] };
  assign truncR_161 = truncval_imm_174;
  wire [28-1:0] truncR_shift_175;
  assign truncR_shift_175 = truncR_161 >>> 94;
  wire [28-1:0] truncR_imm_176;
  assign truncR_imm_176 = (truncR_161[121])? truncR_shift_175[27:0] : truncR_161[121:94];
  assign padl_bits_160 = truncR_imm_176;
  assign padl_159 = { { 5{ padl_bits_160[27] } }, padl_bits_160 };
  assign truncR_158 = padl_159;
  wire [31-1:0] truncR_shift_177;
  assign truncR_shift_177 = truncR_158 >>> 2;
  wire [31-1:0] truncR_imm_178;
  assign truncR_imm_178 = (truncR_158[32])? truncR_shift_177[30:0] : truncR_158[32:2];
  wire [40-1:0] truncR_179;
  wire [40-1:0] padl_180;
  wire [35-1:0] padl_bits_181;
  wire [122-1:0] truncR_182;
  wire [135-1:0] truncval_183;
  wire [135-1:0] padl_184;
  wire [67-1:0] padl_bits_185;
  wire [67-1:0] padl_186;
  wire [61-1:0] padl_bits_187;
  wire [1-1:0] toSInt_188;
  assign toSInt_188 = 0;
  wire [61-1:0] toSInt_imm_189;
  wire [60-1:0] const_190;
  assign const_190 = 60'd57646075230342;
  assign toSInt_imm_189 = { toSInt_188, const_190 };
  assign padl_bits_187 = toSInt_imm_189;
  assign padl_186 = { { 6{ padl_bits_187[60] } }, padl_bits_187 };
  assign padl_bits_185 = padl_186;
  assign padl_184 = { { 68{ padl_bits_185[66] } }, padl_bits_185 };
  wire [135-1:0] padl_191;
  wire [67-1:0] padl_bits_192;
  wire [67-1:0] padr_193;
  wire [41-1:0] padr_bits_194;
  assign padr_bits_194 = 0;
  assign padr_193 = { dxdt, padr_bits_194 };
  assign padl_bits_192 = padr_193;
  assign padl_191 = { { 68{ padl_bits_192[66] } }, padl_bits_192 };
  assign truncval_183 = padl_184 * padl_191;
  wire [122-1:0] truncval_imm_195;
  assign truncval_imm_195 = { truncval_183[134], truncval_183[120:0] };
  assign truncR_182 = truncval_imm_195;
  wire [35-1:0] truncR_shift_196;
  assign truncR_shift_196 = truncR_182 >>> 87;
  wire [35-1:0] truncR_imm_197;
  assign truncR_imm_197 = (truncR_182[121])? truncR_shift_196[34:0] : truncR_182[121:87];
  assign padl_bits_181 = truncR_imm_197;
  assign padl_180 = { { 5{ padl_bits_181[34] } }, padl_bits_181 };
  assign truncR_179 = padl_180;
  wire [31-1:0] truncR_shift_198;
  assign truncR_shift_198 = truncR_179 >>> 9;
  wire [31-1:0] truncR_imm_199;
  assign truncR_imm_199 = (truncR_179[39])? truncR_shift_198[30:0] : truncR_179[39:9];

  always @(posedge clk) begin
    if(reset) begin
      prev_input_voltage_real <= 0;
    end else begin
      prev_input_voltage_real <= input_voltage_real;
    end
    if(reset | (1'd0 | (prev_input_voltage_real - input_voltage_real != 0))) begin
      input_voltage_prev <= 10'd0;
    end else begin
      input_voltage_prev <= input_voltage_real;
    end
    if(reset | (1'd0 | (prev_input_voltage_real - input_voltage_real != 0))) begin
      v <= 31'd0;
    end else begin
      v <= v + truncR_imm_178;
    end
    if(reset | (1'd0 | (prev_input_voltage_real - input_voltage_real != 0))) begin
      x <= 31'd16777216;
    end else begin
      x <= x + truncR_imm_199;
    end
  end


endmodule


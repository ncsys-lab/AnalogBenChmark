

module voltage_controlled_oscillator #
(
  parameter gain = 1536,
  parameter damping_resistance = 1228
)
(
  input clk,
  input reset,
  input [10-1:0] input_voltage_real,
  output [12-1:0] output_clock_real
);

  reg [12-1:0] x;
  reg [12-1:0] v;
  wire [9-1:0] dvdt;
  wire [9-1:0] dxdt;
  wire [19-1:0] truncR_0;
  wire [25-1:0] truncval_1;
  wire [25-1:0] padl_2;
  wire [12-1:0] padl_bits_3;
  wire [12-1:0] padr_4;
  wire [2-1:0] padr_bits_5;
  assign padr_bits_5 = 0;
  wire [10-1:0] neg_imm_6;
  wire [27-1:0] truncR_7;
  wire [35-1:0] truncval_8;
  wire [35-1:0] padl_9;
  wire [17-1:0] padl_bits_10;
  wire [17-1:0] padr_11;
  wire [7-1:0] padr_bits_12;
  assign padr_bits_12 = 0;
  wire [20-1:0] truncR_13;
  wire [21-1:0] truncval_14;
  wire [21-1:0] padl_15;
  wire [10-1:0] padl_bits_16;
  wire [10-1:0] padr_17;
  wire [1-1:0] padr_bits_18;
  assign padr_bits_18 = 0;
  wire [9-1:0] padl_19;
  wire [8-1:0] padl_bits_20;
  wire [24-1:0] truncR_21;
  wire [28-1:0] truncval_22;
  wire [28-1:0] padl_23;
  wire [14-1:0] padl_bits_24;
  wire [14-1:0] padl_25;
  wire [11-1:0] padl_bits_26;
  wire [11-1:0] param_27;
  assign param_27 = gain;
  assign padl_bits_26 = param_27;
  wire [3-1:0] padl_bits_zero_28;
  assign padl_bits_zero_28 = 0;
  assign padl_25 = { padl_bits_zero_28, padl_bits_26 };
  assign padl_bits_24 = padl_25;
  wire [14-1:0] padl_bits_zero_29;
  assign padl_bits_zero_29 = 0;
  assign padl_23 = { padl_bits_zero_29, padl_bits_24 };
  wire [28-1:0] padl_30;
  wire [14-1:0] padl_bits_31;
  wire [14-1:0] padr_32;
  wire [4-1:0] padr_bits_33;
  assign padr_bits_33 = 0;
  assign padr_32 = { input_voltage_real, padr_bits_33 };
  assign padl_bits_31 = padr_32;
  wire [14-1:0] padl_bits_zero_34;
  assign padl_bits_zero_34 = 0;
  assign padl_30 = { padl_bits_zero_34, padl_bits_31 };
  assign truncval_22 = padl_23 * padl_30;
  assign truncR_21 = truncval_22[23:0];
  assign padl_bits_20 = truncR_21[23:16];
  wire [1-1:0] padl_bits_zero_35;
  assign padl_bits_zero_35 = 0;
  assign padl_19 = { padl_bits_zero_35, padl_bits_20 };
  assign padr_17 = { padl_19, padr_bits_18 };
  assign padl_bits_16 = padr_17;
  wire [11-1:0] padl_bits_zero_36;
  assign padl_bits_zero_36 = 0;
  assign padl_15 = { padl_bits_zero_36, padl_bits_16 };
  wire [21-1:0] padl_37;
  wire [10-1:0] padl_bits_38;
  assign padl_bits_38 = input_voltage_real;
  wire [11-1:0] padl_bits_zero_39;
  assign padl_bits_zero_39 = 0;
  assign padl_37 = { padl_bits_zero_39, padl_bits_38 };
  assign truncval_14 = padl_15 * padl_37;
  wire [20-1:0] truncval_imm_40;
  assign truncval_imm_40 = { truncval_14[20], truncval_14[18:0] };
  assign truncR_13 = truncval_imm_40;
  wire [10-1:0] truncR_shift_41;
  assign truncR_shift_41 = truncR_13 >>> 10;
  wire [10-1:0] truncR_imm_42;
  assign truncR_imm_42 = (truncR_13[19])? truncR_shift_41[9:0] : truncR_13[19:10];
  assign padr_11 = { truncR_imm_42, padr_bits_12 };
  assign padl_bits_10 = padr_11;
  assign padl_9 = { { 18{ padl_bits_10[16] } }, padl_bits_10 };
  wire [35-1:0] padl_43;
  wire [17-1:0] padl_bits_44;
  wire [17-1:0] padl_45;
  wire [12-1:0] padl_bits_46;
  wire [1-1:0] toSInt_47;
  assign toSInt_47 = 0;
  wire [12-1:0] toSInt_imm_48;
  wire [11-1:0] param_49;
  assign param_49 = gain;
  assign toSInt_imm_48 = { toSInt_47, param_49 };
  assign padl_bits_46 = toSInt_imm_48;
  assign padl_45 = { { 5{ padl_bits_46[11] } }, padl_bits_46 };
  assign padl_bits_44 = padl_45;
  assign padl_43 = { { 18{ padl_bits_44[16] } }, padl_bits_44 };
  assign truncval_8 = padl_9 * padl_43;
  wire [27-1:0] truncval_imm_50;
  assign truncval_imm_50 = { truncval_8[34], truncval_8[25:0] };
  assign truncR_7 = truncval_imm_50;
  wire [10-1:0] truncR_shift_51;
  assign truncR_shift_51 = truncR_7 >>> 17;
  wire [10-1:0] truncR_imm_52;
  assign truncR_imm_52 = (truncR_7[26])? truncR_shift_51[9:0] : truncR_7[26:17];
  assign neg_imm_6 = -truncR_imm_52;
  assign padr_4 = { neg_imm_6, padr_bits_5 };
  assign padl_bits_3 = padr_4;
  assign padl_2 = { { 13{ padl_bits_3[11] } }, padl_bits_3 };
  wire [25-1:0] padl_53;
  wire [12-1:0] padl_bits_54;
  assign padl_bits_54 = x;
  assign padl_53 = { { 13{ padl_bits_54[11] } }, padl_bits_54 };
  assign truncval_1 = padl_2 * padl_53;
  wire [19-1:0] truncval_imm_55;
  assign truncval_imm_55 = { truncval_1[24], truncval_1[17:0] };
  assign truncR_0 = truncval_imm_55;
  wire [9-1:0] truncR_shift_56;
  assign truncR_shift_56 = truncR_0 >>> 10;
  wire [9-1:0] truncR_imm_57;
  assign truncR_imm_57 = (truncR_0[18])? truncR_shift_56[8:0] : truncR_0[18:10];
  assign dvdt = truncR_imm_57;
  wire [12-1:0] truncR_58;
  assign truncR_58 = v;
  wire [9-1:0] truncR_shift_59;
  assign truncR_shift_59 = truncR_58 >>> 3;
  wire [9-1:0] truncR_imm_60;
  assign truncR_imm_60 = (truncR_58[11])? truncR_shift_59[8:0] : truncR_58[11:3];
  assign dxdt = truncR_imm_60;
  assign output_clock_real = x;
  wire [15-1:0] truncR_61;
  wire [15-1:0] padl_62;
  wire [12-1:0] padl_bits_63;
  wire [40-1:0] truncR_64;
  wire [49-1:0] truncval_65;
  wire [49-1:0] padl_66;
  wire [24-1:0] padl_bits_67;
  wire [24-1:0] padl_68;
  wire [20-1:0] padl_bits_69;
  wire [1-1:0] toSInt_70;
  assign toSInt_70 = 0;
  wire [20-1:0] toSInt_imm_71;
  wire [19-1:0] const_72;
  assign const_72 = 5242;
  assign toSInt_imm_71 = { toSInt_70, const_72 };
  assign padl_bits_69 = toSInt_imm_71;
  assign padl_68 = { { 4{ padl_bits_69[19] } }, padl_bits_69 };
  assign padl_bits_67 = padl_68;
  assign padl_66 = { { 25{ padl_bits_67[23] } }, padl_bits_67 };
  wire [49-1:0] padl_73;
  wire [24-1:0] padl_bits_74;
  wire [24-1:0] padr_75;
  wire [15-1:0] padr_bits_76;
  assign padr_bits_76 = 0;
  assign padr_75 = { dvdt, padr_bits_76 };
  assign padl_bits_74 = padr_75;
  assign padl_73 = { { 25{ padl_bits_74[23] } }, padl_bits_74 };
  assign truncval_65 = padl_66 * padl_73;
  wire [40-1:0] truncval_imm_77;
  assign truncval_imm_77 = { truncval_65[48], truncval_65[38:0] };
  assign truncR_64 = truncval_imm_77;
  wire [12-1:0] truncR_shift_78;
  assign truncR_shift_78 = truncR_64 >>> 28;
  wire [12-1:0] truncR_imm_79;
  assign truncR_imm_79 = (truncR_64[39])? truncR_shift_78[11:0] : truncR_64[39:28];
  assign padl_bits_63 = truncR_imm_79;
  assign padl_62 = { { 3{ padl_bits_63[11] } }, padl_bits_63 };
  assign truncR_61 = padl_62;
  wire [12-1:0] truncR_shift_80;
  assign truncR_shift_80 = truncR_61 >>> 3;
  wire [12-1:0] truncR_imm_81;
  assign truncR_imm_81 = (truncR_61[14])? truncR_shift_80[11:0] : truncR_61[14:3];
  wire [16-1:0] truncR_82;
  wire [16-1:0] padl_83;
  wire [13-1:0] padl_bits_84;
  wire [40-1:0] truncR_85;
  wire [49-1:0] truncval_86;
  wire [49-1:0] padl_87;
  wire [24-1:0] padl_bits_88;
  wire [24-1:0] padl_89;
  wire [20-1:0] padl_bits_90;
  wire [1-1:0] toSInt_91;
  assign toSInt_91 = 0;
  wire [20-1:0] toSInt_imm_92;
  wire [19-1:0] const_93;
  assign const_93 = 5242;
  assign toSInt_imm_92 = { toSInt_91, const_93 };
  assign padl_bits_90 = toSInt_imm_92;
  assign padl_89 = { { 4{ padl_bits_90[19] } }, padl_bits_90 };
  assign padl_bits_88 = padl_89;
  assign padl_87 = { { 25{ padl_bits_88[23] } }, padl_bits_88 };
  wire [49-1:0] padl_94;
  wire [24-1:0] padl_bits_95;
  wire [24-1:0] padr_96;
  wire [13-1:0] padr_bits_97;
  assign padr_bits_97 = 0;
  wire [11-1:0] padr_98;
  wire [2-1:0] padr_bits_99;
  assign padr_bits_99 = 0;
  assign padr_98 = { dxdt, padr_bits_99 };
  wire [11-1:0] padl_100;
  wire [9-1:0] padl_bits_101;
  wire [27-1:0] truncR_102;
  wire [35-1:0] truncval_103;
  wire [35-1:0] padl_104;
  wire [17-1:0] padl_bits_105;
  wire [17-1:0] padl_106;
  wire [13-1:0] padl_bits_107;
  wire [1-1:0] toSInt_108;
  assign toSInt_108 = 0;
  wire [13-1:0] toSInt_imm_109;
  wire [12-1:0] param_110;
  assign param_110 = damping_resistance;
  assign toSInt_imm_109 = { toSInt_108, param_110 };
  assign padl_bits_107 = toSInt_imm_109;
  assign padl_106 = { { 4{ padl_bits_107[12] } }, padl_bits_107 };
  assign padl_bits_105 = padl_106;
  assign padl_104 = { { 18{ padl_bits_105[16] } }, padl_bits_105 };
  wire [35-1:0] padl_111;
  wire [17-1:0] padl_bits_112;
  wire [17-1:0] padr_113;
  wire [5-1:0] padr_bits_114;
  assign padr_bits_114 = 0;
  assign padr_113 = { v, padr_bits_114 };
  assign padl_bits_112 = padr_113;
  assign padl_111 = { { 18{ padl_bits_112[16] } }, padl_bits_112 };
  assign truncval_103 = padl_104 * padl_111;
  wire [27-1:0] truncval_imm_115;
  assign truncval_imm_115 = { truncval_103[34], truncval_103[25:0] };
  assign truncR_102 = truncval_imm_115;
  wire [9-1:0] truncR_shift_116;
  assign truncR_shift_116 = truncR_102 >>> 18;
  wire [9-1:0] truncR_imm_117;
  assign truncR_imm_117 = (truncR_102[26])? truncR_shift_116[8:0] : truncR_102[26:18];
  assign padl_bits_101 = truncR_imm_117;
  assign padl_100 = { { 2{ padl_bits_101[8] } }, padl_bits_101 };
  assign padr_96 = { padr_98 - padl_100, padr_bits_97 };
  assign padl_bits_95 = padr_96;
  assign padl_94 = { { 25{ padl_bits_95[23] } }, padl_bits_95 };
  assign truncval_86 = padl_87 * padl_94;
  wire [40-1:0] truncval_imm_118;
  assign truncval_imm_118 = { truncval_86[48], truncval_86[38:0] };
  assign truncR_85 = truncval_imm_118;
  wire [13-1:0] truncR_shift_119;
  assign truncR_shift_119 = truncR_85 >>> 27;
  wire [13-1:0] truncR_imm_120;
  assign truncR_imm_120 = (truncR_85[39])? truncR_shift_119[12:0] : truncR_85[39:27];
  assign padl_bits_84 = truncR_imm_120;
  assign padl_83 = { { 3{ padl_bits_84[12] } }, padl_bits_84 };
  assign truncR_82 = padl_83;
  wire [12-1:0] truncR_shift_121;
  assign truncR_shift_121 = truncR_82 >>> 4;
  wire [12-1:0] truncR_imm_122;
  assign truncR_imm_122 = (truncR_82[15])? truncR_shift_121[11:0] : truncR_82[15:4];

  always @(posedge clk) begin
    if(reset) begin
      v <= 0;
    end else begin
      v <= v + truncR_imm_81;
    end
    if(reset) begin
      x <= 128;
    end else begin
      x <= x + truncR_imm_122;
    end
  end


endmodule

